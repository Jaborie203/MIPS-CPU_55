`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:34:24 05/06/2016 
// Design Name: 
// Module Name:    decoder5_32 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module decoder5_32(
    input [4:0] data_in,
    input ena,
    output reg[31:0] data_out
    );
    //reg[31:0] data_temp;
    //assign data_out = data_temp;
    always @ (ena or data_in) begin
    if (ena == 1)
	    case(data_in)
		    5'b00000:
                 data_out= 32'b11111111111111111111111111111110;
		    5'b00001:
                 data_out= 32'b11111111111111111111111111111101;
		    5'b00010:
                 data_out= 32'b11111111111111111111111111111011;
		    5'b00011:
                 data_out= 32'b11111111111111111111111111110111;
		    5'b00100:
                 data_out= 32'b11111111111111111111111111101111;
		    5'b00101:
                 data_out= 32'b11111111111111111111111111011111;
		    5'b00110:
                 data_out= 32'b11111111111111111111111110111111;
		    5'b00111:
                 data_out= 32'b11111111111111111111111101111111;
			 5'b01000:
                 data_out= 32'b11111111111111111111111011111111;
		    5'b01001:
                 data_out= 32'b11111111111111111111110111111111;
		    5'b01010:
                 data_out= 32'b11111111111111111111101111111111;
		    5'b01011:
                 data_out= 32'b11111111111111111111011111111111;
		    5'b01100:
                 data_out= 32'b11111111111111111110111111111111;
		    5'b01101:
                 data_out= 32'b11111111111111111101111111111111;
		    5'b01110:
                 data_out= 32'b11111111111111111011111111111111;
		    5'b01111:
                 data_out= 32'b11111111111111110111111111111111;
			 5'b10000:
                 data_out= 32'b11111111111111101111111111111111;
		    5'b10001:
                 data_out= 32'b11111111111111011111111111111111;
		    5'b10010:
                 data_out= 32'b11111111111110111111111111111111;
		    5'b10011:
                 data_out= 32'b11111111111101111111111111111111;
		    5'b10100:
                 data_out= 32'b11111111111011111111111111111111;
		    5'b10101:
                 data_out= 32'b11111111110111111111111111111111;
		    5'b10110:
                 data_out= 32'b11111111101111111111111111111111;
		    5'b10111:
                 data_out= 32'b11111111011111111111111111111111;
			 5'b11000:
                 data_out= 32'b11111110111111111111111111111111;
		    5'b11001:
                 data_out= 32'b11111101111111111111111111111111;
		    5'b11010:
                 data_out= 32'b11111011111111111111111111111111;
		    5'b11011:
                 data_out= 32'b11110111111111111111111111111111;
		    5'b11100:
                 data_out= 32'b11101111111111111111111111111111;
		    5'b11101:
                 data_out= 32'b11011111111111111111111111111111;
		    5'b11110:
                 data_out= 32'b10111111111111111111111111111111;
		    5'b11111:
                 data_out= 32'b01111111111111111111111111111111;
       endcase
    else
       data_out = 32'b11111111111111111111111111111111;
    end
endmodule

