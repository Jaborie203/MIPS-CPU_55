`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:36:30 05/03/2016 
// Design Name: 
// Module Name:    sccomp_dataflow 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module sccomp_dataflow(clock,reset,pc_out,inst,aluout,dmemout);
    input clock,reset;
	 output [31:0] pc_out,inst,aluout,dmemout;
	 wire [31:0] dmemdata;
	 wire dmemwena;
	 wire [1:0]wbh;
	 wire wbh_fh;
	 
	 sccpu_dataflow cpu(clock,reset,pc_out,inst,dmemwena,aluout,dmemdata,dmemout,wbh,wbh_fh);
	 scinstmem imem(pc_out[12:2],inst);
	 scdatamem dmem(clock,wbh,wbh_fh,dmemwena,aluout[12:0],dmemdata,dmemout);//�ڴ�aluout��Ϊ���ݴ洢���ĵ�ַ
endmodule
